* fixed osc subckt
.subckt fixed_osc Out
.include Model_files/2n3904.txt
* DC Power supply
v1 1 0 dc=12
v6 6 0 dc=-12
v11 11 0 dc=-12

* Pitch Tuning signal
vsig5 sig5 0 dc=-2

* Variable Inductor
l6 1 2 94u

c5 1 2 3900p 
c7 2 15 0.01u
c8 1 0 1u 
C6 2 Out 22p
C9 2 8 33p
c10 9 10 1u 
c11 10 0 1u
r9 10 sig5 10k
r10 12 8 470
r11 8 9 33
r12 9 11 10k
r39 10 11 10k
r13 9 0 2.2k
r7 15 5 47k
r8 5 0 1k
r5 4 0 1k
r6 3 6 2.2k

* the BJTs
q1 2 4 3 Q2N3904
q2 1 5 3 Q2N3904
q3 2 12 10 Q2N3904
.ends