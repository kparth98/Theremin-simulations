* detector circuit
.include subvar.cir
.include subfixed.cir
.include Model_files/Diode_1N914.txt

.subckt detector out 
xfixed 1 fixed_osc
xvar 1 var_osc
d1 1 0 1N914
r23 1 out 10k
r24 out 0 47k
c23 out 0 4700p
.ends

* xdetect 1 detector

* .control
* tran 0.1us 5ms
* run

* plot v(1)
* .endc
* .end

