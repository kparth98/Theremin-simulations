.include ina.cir
.include Model_files/ua741.txt
.include detector.cir

vpos dcpos 0 dc = 12
vneg dcneg 0 dc=-12
xina neg pos ref op dcpos dcneg ina
xo 0 2 dcpos dcneg ref ua741

r1 pos sig 180k
r2 neg 0 180k
r3 2 op 10k
c1 ref 2 0.1u

xd sig detector
* vsig sig 0 sin(-3 0.25 2k)

.tran 0.01m 10m
.control
run
plot v(op)
.endc
.end
