detector circuit
.include 2n3904.txt
.include subvar.cir
.include subfixed.cir
.include Diode_1N914.txt
xfixed 3 fixed_osc
xvar 4 var_osc
*v1 3 0 sin(0 5 260k 0 0) dc=1 
*v2 1 0 sin(0 5 260k 0 0) dc=1
*vd1 3 4 dc=0
*vd2 4 1 dc =0
c1 3 1 22p
c2 4 1 22p
d1 1 0 1N914
r23 1 2 10k
r24 2 0 4.7k
c23 2 0 4.7n

.control
tran 0.1us 10us
run
*plotting input and output voltages
plot v(2) 
*v(2)
.endc
.end

