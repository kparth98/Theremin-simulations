test

.include detector.cir

xd 1 detector

.tran 0.1u 1m

.control
run
plot v(1)
.endc
.end