vca processor
.include subvol.cir
.include Model_files/LM13700.txt
.include detector.cir
* .include Model_files/Diode_1N914.txt
.include Model_files/1n4148.txt
.include vca_new.cir

* xd1 16 15 0 13 12 6 10 9 11 LM13600/NS
.subckt vca_proc vol op
xd1 16 15 0 vol op 6 10 9 11 lm13700/ns
v1 6 0 dc=-12
v2 11 0 dc=12
* vvol vol 0 sin(0 10 450k)
r35 11 vol 1.8Meg
r36 11 15 1.8Meg
c27 vol 0 0.1u
r37 vol t 4.7Meg
xd t op 1n4148
r38 11 16 47k
.ends

* xvol vol vol_osc
vvol vol 0 dc=11.3
xproc vol vca_pro vca_proc
*12 goes to VCA 
*10 is the audio output
* v12 12 0 dc=-4
* .subckt vca audio dtc vca_proc
* xd2 1 2 dtc 4 5 6 7 8 11 lm13700/ns
* * * vinp 3 0 sin(0 2 1k) dc=-1
* xdetect 3 detector
* vshort 5 7 dc=0
* r25 4 6 330k
* r26 4 0 4.7k
* r27 2 sig9 100k
* r28 4 sig7 150k
* r29 1 6 100k
* r30 1 vca_proc 47k
* r31	5 0 4.7k
* r32 8 6 4.7k
* c24 7 0 3.3n
* c25 8 t2 1u
* r33 t2 audio 4.7k
* c26 audio 0 0.01u
* r34 audio 0 4.7k
* .ends
xdtc dtc detector
xvca audio dtc vca_pro vca

.control
tran 0.01m 10m
run
* plot v(3) v(10) v(12) v(13)
plot v(audio) 
plot v(dtc) v(vca_pro) v(audio)

.endc
.end
