* subcircuit volume oscillator
.include Model_files/2n3904.txt
* .include Model_files/Diode_1N914.txt
.include Model_files/1n4148.txt

.subckt vol_osc Out
* the volume antenna circuit
la a 1 12.5m
ca a 0 15p
xd1 2 1 1N4148
c12 2 3 1000p 
*ic=1
l7 3 1 2.5m
r14 2 Out 560k
v1 4 0 dc=12
v2 9 0 dc=-12
vsig6 sig6 0 dc=-10
*variable inductor
l11 4 5 68u
c13 4 0 1u
c14 5 3 2200p
r17 3 0 470
c15 3 0 0.01u
q1 4 3 6 q2n3904
q2 5 8 6 q2n3904
r15 8 0 470
r16 6 9 2.2k
c16 5 10 22p
r19 10 11 470
q3 5 11 12 q2n3904
c18 12 0 1u
r40 12 9 10k
r18 12 sig6 2.7k
c17 12 13 1u
r21 13 0 2.2k
r22 13 9 10k
r20 13 10 33
.ends